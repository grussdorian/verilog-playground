module example_ckt (z,x,y);
	input x,y;
	output z;
	assign z = x& y;
endmodule

